`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: GDUT
// Engineer: JF Lee
// 
// Create Date:
// Design Name:
// Module Name: 
// Project Name: 
// Taget Devices: zcu104
// Tool Versions: 2018.3
// Description:
// 
// Dependencies:
// 
// Revision: 
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module PE_array#(
	parameter DATA_WIDTH_I = 8,
	parameter DATA_WIDTH_O = 18
)(
	input wire 							clk,
	input wire 							rst,
	
	// input feature map 4 channel
	input wire [3:0]					en_fm,      // fm: feature map
	input wire [DATA_WIDTH_I*25-1:0]	din_fm_c0,
	input wire [DATA_WIDTH_I*25-1:0]	din_fm_c1,
	input wire [DATA_WIDTH_I*25-1:0]	din_fm_c2,
	input wire [DATA_WIDTH_I*25-1:0]	din_fm_c3,
	// input weight 8 batches
	input wire [7:0]					en_w,
	input wire [DATA_WIDTH_I*25-1:0]	din_w_b0,
	input wire [DATA_WIDTH_I*25-1:0]  	din_w_b1,
	input wire [DATA_WIDTH_I*25-1:0]  	din_w_b2,
	input wire [DATA_WIDTH_I*25-1:0]  	din_w_b3,
	input wire [DATA_WIDTH_I*25-1:0]  	din_w_b4,
	input wire [DATA_WIDTH_I*25-1:0]  	din_w_b5,
	input wire [DATA_WIDTH_I*25-1:0]  	din_w_b6,
	input wire [DATA_WIDTH_I*25-1:0]  	din_w_b7,
	
	// output partial sum 0
	output wire	[15:0]					en_psum0,
	output wire [DATA_WIDTH_O*25-1:0]   psum0_pe00,psum0_pe01,psum0_pe02,psum0_pe03,
	output wire [DATA_WIDTH_O*25-1:0]   psum0_pe10,psum0_pe11,psum0_pe12,psum0_pe13,
	output wire [DATA_WIDTH_O*25-1:0]   psum0_pe20,psum0_pe21,psum0_pe22,psum0_pe23,
	output wire [DATA_WIDTH_O*25-1:0]   psum0_pe30,psum0_pe31,psum0_pe32,psum0_pe33,
	// output partial sum 1
	output wire	[15:0]					en_psum1,
	output wire [DATA_WIDTH_O*25-1:0]   psum1_pe00,psum1_pe01,psum1_pe02,psum1_pe03,
	output wire [DATA_WIDTH_O*25-1:0]   psum1_pe10,psum1_pe11,psum1_pe12,psum1_pe13,
	output wire [DATA_WIDTH_O*25-1:0]   psum1_pe20,psum1_pe21,psum1_pe22,psum1_pe23,
	output wire [DATA_WIDTH_O*25-1:0]   psum1_pe30,psum1_pe31,psum1_pe32,psum1_pe33
);
	wire						en_out_fm_pe00,en_out_fm_pe01,en_out_fm_pe02;
	wire						en_out_fm_pe10,en_out_fm_pe11,en_out_fm_pe12;
	wire						en_out_fm_pe20,en_out_fm_pe21,en_out_fm_pe22;
	wire						en_out_fm_pe30,en_out_fm_pe31,en_out_fm_pe32;
	
	wire						en_out_w_b0_pe00,en_out_w_b0_pe01,en_out_w_b0_pe02,en_out_w_b0_pe03;
	wire						en_out_w_b0_pe10,en_out_w_b0_pe11,en_out_w_b0_pe12,en_out_w_b0_pe13;
	wire						en_out_w_b0_pe20,en_out_w_b0_pe21,en_out_w_b0_pe22,en_out_w_b0_pe23;
	
	wire						en_out_w_b1_pe00,en_out_w_b1_pe01,en_out_w_b1_pe02,en_out_w_b1_pe03;
	wire						en_out_w_b1_pe10,en_out_w_b1_pe11,en_out_w_b1_pe12,en_out_w_b1_pe13;
	wire						en_out_w_b1_pe20,en_out_w_b1_pe21,en_out_w_b1_pe22,en_out_w_b1_pe23;
	
	wire [DATA_WIDTH_I*25-1:0]	dout_fm_pe00,dout_fm_pe01,dout_fm_pe02;
	wire [DATA_WIDTH_I*25-1:0]	dout_fm_pe10,dout_fm_pe11,dout_fm_pe12;
	wire [DATA_WIDTH_I*25-1:0]	dout_fm_pe20,dout_fm_pe21,dout_fm_pe22;
	wire [DATA_WIDTH_I*25-1:0]	dout_fm_pe30,dout_fm_pe31,dout_fm_pe32;
	
	wire [DATA_WIDTH_I*25-1:0]	dout_w_b0_pe00,dout_w_b0_pe01,dout_w_b0_pe02,dout_w_b0_pe03;
	wire [DATA_WIDTH_I*25-1:0]	dout_w_b0_pe10,dout_w_b0_pe11,dout_w_b0_pe12,dout_w_b0_pe13;
	wire [DATA_WIDTH_I*25-1:0]	dout_w_b0_pe20,dout_w_b0_pe21,dout_w_b0_pe22,dout_w_b0_pe23;
	
	wire [DATA_WIDTH_I*25-1:0]	dout_w_b1_pe00,dout_w_b1_pe01,dout_w_b1_pe02,dout_w_b1_pe03;
	wire [DATA_WIDTH_I*25-1:0]	dout_w_b1_pe10,dout_w_b1_pe11,dout_w_b1_pe12,dout_w_b1_pe13;
	wire [DATA_WIDTH_I*25-1:0]	dout_w_b1_pe20,dout_w_b1_pe21,dout_w_b1_pe22,dout_w_b1_pe23;

	(* keep = "true" *)
	reg rst_d1;
	always@(posedge clk)begin
		if(rst)begin
			rst_d1 <= 1'b1;
		end
		else begin
			rst_d1 <= 1'b0;
		end
	end

pe_norm#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
)pe_00(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_fm[0]), // ok
	.din_fm_00(din_fm_c0[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(din_fm_c0[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(din_fm_c0[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(din_fm_c0[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(din_fm_c0[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(din_fm_c0[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(din_fm_c0[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(din_fm_c0[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(din_fm_c0[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(din_fm_c0[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(din_fm_c0[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(din_fm_c0[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(din_fm_c0[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(din_fm_c0[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(din_fm_c0[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(din_fm_c0[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(din_fm_c0[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_fm_32(din_fm_c0[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(din_fm_c0[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(din_fm_c0[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(din_fm_c0[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(din_fm_c0[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(din_fm_c0[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(din_fm_c0[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(din_fm_c0[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_w[0]), // ok
	.din_w_b0_00(din_w_b0[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(din_w_b0[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(din_w_b0[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(din_w_b0[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(din_w_b0[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(din_w_b0[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(din_w_b0[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(din_w_b0[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(din_w_b0[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(din_w_b0[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(din_w_b0[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(din_w_b0[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(din_w_b0[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(din_w_b0[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(din_w_b0[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(din_w_b0[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(din_w_b0[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b0_32(din_w_b0[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(din_w_b0[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(din_w_b0[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(din_w_b0[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(din_w_b0[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(din_w_b0[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(din_w_b0[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(din_w_b0[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_w[4]), // ok
	.din_w_b1_00(din_w_b1[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(din_w_b1[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(din_w_b1[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(din_w_b1[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(din_w_b1[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(din_w_b1[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(din_w_b1[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(din_w_b1[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(din_w_b1[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(din_w_b1[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(din_w_b1[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(din_w_b1[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(din_w_b1[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(din_w_b1[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(din_w_b1[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(din_w_b1[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(din_w_b1[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(din_w_b1[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(din_w_b1[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(din_w_b1[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(din_w_b1[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(din_w_b1[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(din_w_b1[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(din_w_b1[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(din_w_b1[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe00), // ok
	.dout_fm_00(dout_fm_pe00[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe00[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe00[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe00[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe00[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe00[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe00[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe00[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe00[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe00[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe00[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe00[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe00[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe00[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe00[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe00[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe00[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe00[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe00[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe00[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe00[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe00[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe00[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe00[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe00[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe00), // ok
	.dout_w_b0_00(dout_w_b0_pe00[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe00[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe00[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe00[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_w_b0_04(dout_w_b0_pe00[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe00[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe00[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe00[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe00[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe00[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe00[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe00[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe00[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe00[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe00[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe00[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe00[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe00[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe00[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe00[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe00[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe00[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe00[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe00[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b0_44(dout_w_b0_pe00[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk
	.en_out_w_b1(en_out_w_b1_pe00), // ok
	.dout_w_b1_00(dout_w_b1_pe00[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe00[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe00[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe00[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_w_b1_04(dout_w_b1_pe00[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe00[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe00[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe00[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe00[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe00[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe00[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe00[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe00[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe00[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe00[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b1_30(dout_w_b1_pe00[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe00[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe00[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe00[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe00[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe00[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe00[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe00[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe00[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe00[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0
	.en_psum0(en_psum0[0]), // ok
	.dout_psum0_00(psum0_pe00[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe00[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe00[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe00[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe00[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe00[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe00[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe00[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe00[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe00[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum0_20(psum0_pe00[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe00[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum0_22(psum0_pe00[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe00[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe00[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),
	.dout_psum0_30(psum0_pe00[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe00[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe00[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe00[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe00[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),
	.dout_psum0_40(psum0_pe00[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe00[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe00[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe00[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe00[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1
	.en_psum1(en_psum1[0]), // ok
	.dout_psum1_00(psum1_pe00[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe00[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe00[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe00[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe00[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe00[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe00[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe00[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe00[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe00[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe00[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe00[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe00[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe00[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe00[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),
	.dout_psum1_30(psum1_pe00[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe00[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe00[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe00[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe00[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),
	.dout_psum1_40(psum1_pe00[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe00[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe00[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe00[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe00[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_norm#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_01(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe00), // ok
	.din_fm_00(dout_fm_pe00[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe00[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe00[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe00[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe00[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe00[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe00[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe00[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe00[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe00[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe00[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe00[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe00[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe00[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(dout_fm_pe00[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(dout_fm_pe00[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe00[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_fm_32(dout_fm_pe00[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe00[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe00[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe00[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe00[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe00[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe00[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe00[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_w[1]),
	.din_w_b0_00(din_w_b2[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(din_w_b2[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(din_w_b2[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(din_w_b2[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(din_w_b2[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(din_w_b2[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(din_w_b2[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(din_w_b2[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(din_w_b2[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(din_w_b2[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(din_w_b2[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(din_w_b2[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(din_w_b2[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(din_w_b2[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(din_w_b2[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(din_w_b2[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(din_w_b2[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b0_32(din_w_b2[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(din_w_b2[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(din_w_b2[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(din_w_b2[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(din_w_b2[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(din_w_b2[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(din_w_b2[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(din_w_b2[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_w[5]),
	.din_w_b1_00(din_w_b3[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(din_w_b3[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(din_w_b3[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(din_w_b3[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(din_w_b3[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(din_w_b3[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(din_w_b3[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(din_w_b3[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(din_w_b3[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(din_w_b3[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(din_w_b3[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(din_w_b3[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(din_w_b3[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(din_w_b3[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(din_w_b3[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(din_w_b3[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(din_w_b3[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(din_w_b3[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(din_w_b3[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(din_w_b3[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(din_w_b3[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(din_w_b3[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(din_w_b3[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(din_w_b3[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(din_w_b3[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe01),
	.dout_fm_00(dout_fm_pe01[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe01[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe01[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe01[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe01[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe01[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe01[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe01[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe01[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe01[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe01[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe01[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe01[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe01[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe01[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe01[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe01[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe01[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe01[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe01[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe01[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe01[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe01[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe01[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe01[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe01),
	.dout_w_b0_00(dout_w_b0_pe01[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe01[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe01[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe01[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_w_b0_04(dout_w_b0_pe01[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe01[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe01[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe01[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe01[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe01[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe01[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe01[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe01[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe01[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe01[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe01[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe01[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe01[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe01[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe01[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe01[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe01[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe01[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe01[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b0_44(dout_w_b0_pe01[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk
	.en_out_w_b1(en_out_w_b1_pe01),
	.dout_w_b1_00(dout_w_b1_pe01[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe01[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe01[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe01[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_w_b1_04(dout_w_b1_pe01[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe01[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe01[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe01[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe01[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe01[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe01[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe01[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe01[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe01[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe01[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b1_30(dout_w_b1_pe01[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe01[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe01[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe01[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe01[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe01[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe01[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe01[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe01[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe01[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0
	.en_psum0(en_psum0[1]),
	.dout_psum0_00(psum0_pe01[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe01[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe01[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe01[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe01[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe01[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe01[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe01[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe01[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe01[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum0_20(psum0_pe01[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe01[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum0_22(psum0_pe01[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe01[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe01[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe01[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe01[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe01[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe01[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe01[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),
	.dout_psum0_40(psum0_pe01[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe01[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe01[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe01[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe01[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1
	.en_psum1(en_psum1[1]),
	.dout_psum1_00(psum1_pe01[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe01[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe01[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe01[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe01[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe01[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe01[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe01[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe01[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe01[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe01[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe01[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe01[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe01[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe01[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),
	.dout_psum1_30(psum1_pe01[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe01[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe01[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe01[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe01[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),
	.dout_psum1_40(psum1_pe01[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe01[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe01[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe01[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe01[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_norm#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_02(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe01), // ok
	.din_fm_00(dout_fm_pe01[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe01[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe01[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe01[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe01[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe01[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe01[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe01[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe01[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe01[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe01[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe01[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe01[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe01[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),	
	.din_fm_24(dout_fm_pe01[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),	
	.din_fm_30(dout_fm_pe01[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe01[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_fm_32(dout_fm_pe01[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe01[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe01[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe01[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe01[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe01[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe01[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe01[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_w[2]),
	.din_w_b0_00(din_w_b4[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(din_w_b4[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(din_w_b4[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(din_w_b4[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(din_w_b4[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(din_w_b4[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(din_w_b4[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(din_w_b4[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(din_w_b4[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(din_w_b4[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(din_w_b4[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(din_w_b4[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(din_w_b4[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(din_w_b4[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(din_w_b4[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(din_w_b4[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(din_w_b4[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(din_w_b4[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(din_w_b4[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(din_w_b4[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(din_w_b4[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(din_w_b4[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(din_w_b4[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(din_w_b4[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(din_w_b4[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_w[6]),
	.din_w_b1_00(din_w_b5[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(din_w_b5[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(din_w_b5[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(din_w_b5[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(din_w_b5[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(din_w_b5[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(din_w_b5[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(din_w_b5[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(din_w_b5[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(din_w_b5[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(din_w_b5[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(din_w_b5[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(din_w_b5[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(din_w_b5[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(din_w_b5[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(din_w_b5[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(din_w_b5[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(din_w_b5[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(din_w_b5[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(din_w_b5[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(din_w_b5[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(din_w_b5[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(din_w_b5[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(din_w_b5[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(din_w_b5[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe02),
	.dout_fm_00(dout_fm_pe02[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe02[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe02[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe02[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe02[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe02[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe02[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe02[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe02[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe02[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe02[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe02[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe02[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe02[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe02[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe02[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe02[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe02[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe02[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe02[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe02[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe02[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe02[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe02[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe02[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe02),
	.dout_w_b0_00(dout_w_b0_pe02[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe02[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe02[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe02[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_w_b0_04(dout_w_b0_pe02[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe02[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe02[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe02[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe02[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe02[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe02[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe02[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe02[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe02[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe02[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe02[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe02[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe02[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe02[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe02[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe02[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe02[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe02[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe02[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b0_44(dout_w_b0_pe02[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk
	.en_out_w_b1(en_out_w_b1_pe02),
	.dout_w_b1_00(dout_w_b1_pe02[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe02[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe02[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe02[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_w_b1_04(dout_w_b1_pe02[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe02[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe02[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe02[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe02[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe02[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe02[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe02[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe02[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe02[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe02[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b1_30(dout_w_b1_pe02[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe02[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe02[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe02[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe02[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe02[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe02[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe02[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe02[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe02[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0
	.en_psum0(en_psum0[2]),
	.dout_psum0_00(psum0_pe02[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe02[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe02[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe02[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe02[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe02[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe02[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe02[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe02[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe02[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum0_20(psum0_pe02[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe02[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum0_22(psum0_pe02[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe02[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe02[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe02[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe02[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe02[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe02[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe02[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),
	.dout_psum0_40(psum0_pe02[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe02[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe02[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe02[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe02[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1
	.en_psum1(en_psum1[2]),
	.dout_psum1_00(psum1_pe02[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe02[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe02[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe02[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe02[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe02[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe02[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe02[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe02[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe02[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe02[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe02[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe02[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe02[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe02[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),
	.dout_psum1_30(psum1_pe02[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe02[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe02[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe02[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe02[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),
	.dout_psum1_40(psum1_pe02[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe02[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe02[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe02[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe02[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_right#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_03(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe02), // ok
	.din_fm_00(dout_fm_pe02[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe02[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe02[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe02[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe02[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe02[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe02[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe02[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe02[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe02[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe02[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe02[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe02[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe02[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),	
	.din_fm_24(dout_fm_pe02[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),	
	.din_fm_30(dout_fm_pe02[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe02[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_fm_32(dout_fm_pe02[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe02[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe02[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe02[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe02[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe02[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe02[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe02[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_w[3]),
	.din_w_b0_00(din_w_b6[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(din_w_b6[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(din_w_b6[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(din_w_b6[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(din_w_b6[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(din_w_b6[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(din_w_b6[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(din_w_b6[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(din_w_b6[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(din_w_b6[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(din_w_b6[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(din_w_b6[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(din_w_b6[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(din_w_b6[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(din_w_b6[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(din_w_b6[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(din_w_b6[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(din_w_b6[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(din_w_b6[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(din_w_b6[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(din_w_b6[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(din_w_b6[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(din_w_b6[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(din_w_b6[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(din_w_b6[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_w[7]),
	.din_w_b1_00(din_w_b7[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(din_w_b7[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(din_w_b7[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(din_w_b7[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(din_w_b7[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(din_w_b7[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(din_w_b7[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(din_w_b7[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(din_w_b7[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(din_w_b7[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(din_w_b7[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(din_w_b7[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(din_w_b7[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(din_w_b7[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(din_w_b7[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(din_w_b7[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(din_w_b7[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(din_w_b7[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(din_w_b7[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(din_w_b7[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(din_w_b7[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(din_w_b7[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(din_w_b7[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(din_w_b7[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(din_w_b7[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe03),
	.dout_w_b0_00(dout_w_b0_pe03[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe03[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe03[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe03[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_w_b0_04(dout_w_b0_pe03[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe03[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe03[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe03[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe03[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe03[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe03[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe03[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe03[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe03[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe03[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe03[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe03[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe03[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe03[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe03[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe03[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe03[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe03[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe03[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b0_44(dout_w_b0_pe03[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk
	.en_out_w_b1(en_out_w_b1_pe03),
	.dout_w_b1_00(dout_w_b1_pe03[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe03[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe03[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe03[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_w_b1_04(dout_w_b1_pe03[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe03[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe03[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe03[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe03[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe03[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe03[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe03[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe03[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe03[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe03[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b1_30(dout_w_b1_pe03[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe03[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe03[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe03[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe03[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe03[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe03[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe03[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe03[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe03[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0
	.en_psum0(en_psum0[3]),
	.dout_psum0_00(psum0_pe03[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe03[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe03[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe03[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe03[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe03[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe03[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe03[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe03[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe03[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum0_20(psum0_pe03[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe03[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum0_22(psum0_pe03[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe03[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe03[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe03[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe03[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe03[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe03[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe03[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),
	.dout_psum0_40(psum0_pe03[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe03[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe03[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe03[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe03[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1
	.en_psum1(en_psum1[3]),
	.dout_psum1_00(psum1_pe03[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe03[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe03[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe03[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe03[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe03[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe03[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe03[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe03[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe03[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe03[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe03[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe03[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe03[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe03[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),
	.dout_psum1_30(psum1_pe03[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe03[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe03[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe03[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe03[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),
	.dout_psum1_40(psum1_pe03[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe03[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe03[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe03[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe03[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);


pe_norm#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_10(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_fm[1]), // ok
	.din_fm_00(din_fm_c1[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(din_fm_c1[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(din_fm_c1[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(din_fm_c1[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(din_fm_c1[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(din_fm_c1[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(din_fm_c1[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(din_fm_c1[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(din_fm_c1[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(din_fm_c1[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(din_fm_c1[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(din_fm_c1[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(din_fm_c1[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(din_fm_c1[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(din_fm_c1[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(din_fm_c1[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(din_fm_c1[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_fm_32(din_fm_c1[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(din_fm_c1[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(din_fm_c1[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(din_fm_c1[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(din_fm_c1[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(din_fm_c1[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(din_fm_c1[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(din_fm_c1[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe00), // ok
	.din_w_b0_00(dout_w_b0_pe00[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe00[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe00[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe00[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe00[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe00[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe00[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe00[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe00[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe00[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe00[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe00[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe00[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe00[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe00[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe00[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe00[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe00[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe00[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe00[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe00[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe00[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe00[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe00[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe00[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe00), // ok
	.din_w_b1_00(dout_w_b1_pe00[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe00[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe00[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe00[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe00[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe00[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe00[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe00[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe00[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe00[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe00[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe00[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe00[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe00[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe00[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe00[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe00[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe00[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe00[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe00[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe00[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe00[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe00[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe00[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe00[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe10),
	.dout_fm_00(dout_fm_pe10[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe10[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe10[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe10[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe10[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe10[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe10[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe10[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe10[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe10[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe10[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe10[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe10[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe10[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe10[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe10[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe10[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe10[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe10[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe10[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe10[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe10[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe10[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe10[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe10[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe10),
	.dout_w_b0_00(dout_w_b0_pe10[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe10[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe10[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe10[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b0_04(dout_w_b0_pe10[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe10[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe10[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe10[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe10[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe10[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe10[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe10[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe10[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe10[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe10[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe10[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe10[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe10[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe10[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe10[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe10[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe10[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe10[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe10[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),	
	.dout_w_b0_44(dout_w_b0_pe10[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk	
	.en_out_w_b1(en_out_w_b1_pe10),
	.dout_w_b1_00(dout_w_b1_pe10[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe10[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe10[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe10[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b1_04(dout_w_b1_pe10[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe10[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe10[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe10[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe10[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe10[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe10[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe10[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe10[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe10[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe10[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),	
	.dout_w_b1_30(dout_w_b1_pe10[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe10[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe10[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe10[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe10[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe10[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe10[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe10[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe10[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe10[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[4]),
	.dout_psum0_00(psum0_pe10[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe10[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe10[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe10[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe10[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe10[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe10[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe10[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe10[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe10[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe10[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe10[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe10[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe10[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe10[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe10[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe10[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe10[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe10[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe10[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe10[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe10[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe10[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe10[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe10[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[4]),
	.dout_psum1_00(psum1_pe10[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe10[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe10[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe10[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe10[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe10[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe10[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe10[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe10[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe10[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe10[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe10[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe10[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe10[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe10[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe10[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe10[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe10[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe10[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe10[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe10[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe10[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe10[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe10[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe10[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_norm#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_11(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe10),
	.din_fm_00(dout_fm_pe10[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe10[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe10[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe10[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe10[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe10[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe10[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe10[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe10[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe10[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe10[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe10[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe10[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe10[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(dout_fm_pe10[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(dout_fm_pe10[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe10[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_fm_32(dout_fm_pe10[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe10[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe10[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe10[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe10[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe10[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe10[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe10[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe01),
	.din_w_b0_00(dout_w_b0_pe01[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe01[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe01[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe01[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe01[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe01[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe01[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe01[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe01[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe01[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe01[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe01[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe01[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe01[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe01[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe01[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe01[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe01[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe01[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe01[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe01[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe01[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe01[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe01[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe01[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe01),
	.din_w_b1_00(dout_w_b1_pe01[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe01[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe01[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe01[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe01[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe01[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe01[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe01[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe01[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe01[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe01[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe01[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe01[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe01[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe01[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe01[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe01[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe01[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe01[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe01[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe01[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe01[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe01[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe01[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe01[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe11),
	.dout_fm_00(dout_fm_pe11[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe11[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe11[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe11[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe11[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe11[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe11[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe11[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe11[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe11[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe11[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe11[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe11[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe11[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe11[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe11[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe11[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe11[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe11[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe11[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe11[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe11[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe11[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe11[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe11[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe11),
	.dout_w_b0_00(dout_w_b0_pe11[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe11[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe11[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe11[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b0_04(dout_w_b0_pe11[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe11[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe11[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe11[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe11[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe11[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe11[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe11[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe11[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe11[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe11[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe11[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe11[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe11[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe11[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe11[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe11[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe11[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe11[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe11[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),	
	.dout_w_b0_44(dout_w_b0_pe11[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk	
	.en_out_w_b1(en_out_w_b1_pe11),
	.dout_w_b1_00(dout_w_b1_pe11[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe11[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe11[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe11[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b1_04(dout_w_b1_pe11[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe11[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe11[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe11[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe11[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe11[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe11[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe11[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe11[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe11[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe11[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),	
	.dout_w_b1_30(dout_w_b1_pe11[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe11[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe11[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe11[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe11[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe11[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe11[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe11[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe11[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe11[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[5]),
	.dout_psum0_00(psum0_pe11[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe11[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe11[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe11[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe11[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe11[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe11[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe11[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe11[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe11[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe11[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe11[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe11[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe11[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe11[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe11[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe11[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe11[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe11[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe11[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe11[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe11[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe11[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe11[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe11[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[5]),
	.dout_psum1_00(psum1_pe11[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe11[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe11[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe11[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe11[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe11[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe11[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe11[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe11[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe11[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe11[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe11[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe11[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe11[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe11[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe11[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe11[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe11[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe11[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe11[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe11[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe11[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe11[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe11[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe11[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_norm#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_12(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe11),
	.din_fm_00(dout_fm_pe11[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe11[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe11[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe11[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe11[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe11[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe11[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe11[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe11[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe11[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe11[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe11[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe11[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe11[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(dout_fm_pe11[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(dout_fm_pe11[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe11[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_fm_32(dout_fm_pe11[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe11[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe11[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe11[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe11[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe11[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe11[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe11[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe02),
	.din_w_b0_00(dout_w_b0_pe02[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe02[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe02[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe02[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe02[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe02[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe02[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe02[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe02[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe02[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe02[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe02[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe02[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe02[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe02[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe02[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe02[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe02[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe02[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe02[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe02[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe02[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe02[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe02[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe02[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe02),
	.din_w_b1_00(dout_w_b1_pe02[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe02[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe02[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe02[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe02[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe02[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe02[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe02[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe02[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe02[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe02[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe02[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe02[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe02[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe02[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe02[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe02[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe02[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe02[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe02[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe02[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe02[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe02[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe02[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe02[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe12),
	.dout_fm_00(dout_fm_pe12[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe12[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe12[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe12[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe12[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe12[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe12[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe12[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe12[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe12[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe12[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe12[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe12[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe12[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe12[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe12[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe12[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe12[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe12[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe12[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe12[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe12[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe12[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe12[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe12[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe12),
	.dout_w_b0_00(dout_w_b0_pe12[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe12[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe12[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe12[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b0_04(dout_w_b0_pe12[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe12[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe12[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe12[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe12[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe12[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe12[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe12[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe12[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe12[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe12[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe12[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe12[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe12[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe12[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe12[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe12[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe12[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe12[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe12[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),	
	.dout_w_b0_44(dout_w_b0_pe12[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk	
	.en_out_w_b1(en_out_w_b1_pe12),
	.dout_w_b1_00(dout_w_b1_pe12[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe12[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe12[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe12[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b1_04(dout_w_b1_pe12[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe12[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe12[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe12[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe12[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe12[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe12[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe12[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe12[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe12[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe12[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),	
	.dout_w_b1_30(dout_w_b1_pe12[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe12[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe12[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe12[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe12[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe12[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe12[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe12[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe12[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe12[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[6]),
	.dout_psum0_00(psum0_pe12[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe12[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe12[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe12[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe12[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe12[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe12[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe12[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe12[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe12[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe12[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe12[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe12[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe12[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe12[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe12[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe12[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe12[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe12[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe12[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe12[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe12[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe12[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe12[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe12[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[6]),
	.dout_psum1_00(psum1_pe12[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe12[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe12[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe12[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe12[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe12[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe12[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe12[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe12[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe12[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe12[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe12[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe12[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe12[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe12[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe12[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe12[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe12[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe12[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe12[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe12[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe12[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe12[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe12[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe12[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_right#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_13(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe12),
	.din_fm_00(dout_fm_pe12[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe12[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe12[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe12[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe12[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe12[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe12[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe12[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe12[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe12[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe12[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe12[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe12[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe12[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(dout_fm_pe12[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(dout_fm_pe12[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe12[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_fm_32(dout_fm_pe12[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe12[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe12[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe12[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe12[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe12[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe12[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe12[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe03),
	.din_w_b0_00(dout_w_b0_pe03[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe03[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe03[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe03[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe03[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe03[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe03[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe03[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe03[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe03[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe03[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe03[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe03[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe03[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe03[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe03[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe03[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe03[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe03[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe03[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe03[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe03[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe03[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe03[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe03[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe03),
	.din_w_b1_00(dout_w_b1_pe03[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe03[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe03[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe03[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe03[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe03[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe03[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe03[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe03[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe03[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe03[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe03[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe03[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe03[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe03[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe03[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe03[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe03[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe03[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe03[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe03[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe03[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe03[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe03[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe03[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe13),
	.dout_w_b0_00(dout_w_b0_pe13[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe13[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe13[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe13[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b0_04(dout_w_b0_pe13[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe13[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe13[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe13[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe13[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe13[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe13[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe13[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe13[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe13[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe13[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe13[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe13[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe13[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe13[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe13[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe13[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe13[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe13[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe13[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),	
	.dout_w_b0_44(dout_w_b0_pe13[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk	
	.en_out_w_b1(en_out_w_b1_pe13),
	.dout_w_b1_00(dout_w_b1_pe13[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe13[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe13[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe13[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b1_04(dout_w_b1_pe13[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe13[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe13[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe13[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe13[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe13[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe13[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe13[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe13[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe13[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe13[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),	
	.dout_w_b1_30(dout_w_b1_pe13[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe13[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe13[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe13[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe13[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe13[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe13[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe13[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe13[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe13[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[7]),
	.dout_psum0_00(psum0_pe13[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe13[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe13[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe13[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe13[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe13[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe13[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe13[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe13[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe13[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe13[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe13[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe13[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe13[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe13[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe13[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe13[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe13[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe13[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe13[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe13[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe13[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe13[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe13[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe13[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[7]),
	.dout_psum1_00(psum1_pe13[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe13[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe13[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe13[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe13[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe13[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe13[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe13[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe13[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe13[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe13[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe13[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe13[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe13[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe13[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe13[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe13[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe13[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe13[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe13[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe13[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe13[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe13[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe13[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe13[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);


pe_norm#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_20(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_fm[2]),
	.din_fm_00(din_fm_c2[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(din_fm_c2[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(din_fm_c2[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(din_fm_c2[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(din_fm_c2[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(din_fm_c2[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(din_fm_c2[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(din_fm_c2[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(din_fm_c2[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(din_fm_c2[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(din_fm_c2[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(din_fm_c2[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(din_fm_c2[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(din_fm_c2[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(din_fm_c2[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(din_fm_c2[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(din_fm_c2[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_fm_32(din_fm_c2[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(din_fm_c2[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(din_fm_c2[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(din_fm_c2[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(din_fm_c2[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(din_fm_c2[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(din_fm_c2[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(din_fm_c2[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe10),
	.din_w_b0_00(dout_w_b0_pe10[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe10[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe10[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe10[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe10[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe10[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe10[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe10[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe10[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe10[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe10[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe10[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe10[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe10[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe10[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe10[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe10[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe10[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe10[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe10[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe10[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe10[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe10[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe10[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe10[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe10), // ok
	.din_w_b1_00(dout_w_b1_pe10[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe10[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe10[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe10[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe10[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe10[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe10[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe10[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe10[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe10[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe10[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe10[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe10[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe10[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe10[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe10[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe10[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe10[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe10[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe10[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe10[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe10[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe10[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe10[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe10[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe20),
	.dout_fm_00(dout_fm_pe20[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe20[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe20[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe20[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe20[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe20[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe20[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe20[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe20[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe20[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe20[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe20[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe20[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe20[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe20[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe20[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe20[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe20[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe20[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe20[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe20[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe20[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe20[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe20[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe20[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe20),
	.dout_w_b0_00(dout_w_b0_pe20[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe20[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe20[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe20[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b0_04(dout_w_b0_pe20[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe20[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe20[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe20[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe20[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe20[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe20[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe20[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe20[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe20[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe20[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe20[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe20[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe20[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe20[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe20[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe20[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe20[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe20[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe20[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),	
	.dout_w_b0_44(dout_w_b0_pe20[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk	
	.en_out_w_b1(en_out_w_b1_pe20),
	.dout_w_b1_00(dout_w_b1_pe20[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe20[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe20[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe20[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b1_04(dout_w_b1_pe20[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe20[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe20[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe20[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe20[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe20[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe20[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe20[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe20[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe20[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe20[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),	
	.dout_w_b1_30(dout_w_b1_pe20[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe20[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe20[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe20[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe20[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe20[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe20[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe20[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe20[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe20[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[8]),
	.dout_psum0_00(psum0_pe20[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe20[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe20[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe20[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe20[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe20[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe20[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe20[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe20[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe20[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe20[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe20[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe20[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe20[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe20[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe20[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe20[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe20[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe20[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe20[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe20[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe20[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe20[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe20[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe20[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[8]),
	.dout_psum1_00(psum1_pe20[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe20[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe20[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe20[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe20[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe20[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe20[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe20[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe20[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe20[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe20[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe20[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe20[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe20[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe20[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe20[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe20[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe20[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe20[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe20[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe20[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe20[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe20[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe20[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe20[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_norm#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_21(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe20),
	.din_fm_00(dout_fm_pe20[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe20[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe20[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe20[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe20[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe20[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe20[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe20[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe20[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe20[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe20[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe20[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe20[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe20[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(dout_fm_pe20[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(dout_fm_pe20[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe20[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_fm_32(dout_fm_pe20[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe20[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe20[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe20[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe20[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe20[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe20[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe20[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe11),
	.din_w_b0_00(dout_w_b0_pe11[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe11[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe11[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe11[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe11[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe11[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe11[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe11[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe11[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe11[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe11[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe11[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe11[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe11[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe11[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe11[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe11[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe11[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe11[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe11[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe11[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe11[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe11[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe11[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe11[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe11),
	.din_w_b1_00(dout_w_b1_pe11[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe11[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe11[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe11[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe11[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe11[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe11[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe11[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe11[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe11[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe11[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe11[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe11[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe11[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe11[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe11[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe11[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe11[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe11[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe11[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe11[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe11[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe11[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe11[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe11[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe21),
	.dout_fm_00(dout_fm_pe21[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe21[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe21[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe21[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe21[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe21[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe21[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe21[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe21[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe21[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe21[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe21[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe21[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe21[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe21[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe21[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe21[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe21[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe21[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe21[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe21[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe21[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe21[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe21[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe21[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe21),
	.dout_w_b0_00(dout_w_b0_pe21[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe21[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe21[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe21[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b0_04(dout_w_b0_pe21[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe21[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe21[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe21[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe21[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe21[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe21[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe21[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe21[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe21[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe21[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe21[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe21[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe21[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe21[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe21[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe21[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe21[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe21[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe21[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),	
	.dout_w_b0_44(dout_w_b0_pe21[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk	
	.en_out_w_b1(en_out_w_b1_pe21),
	.dout_w_b1_00(dout_w_b1_pe21[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe21[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe21[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe21[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b1_04(dout_w_b1_pe21[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe21[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe21[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe21[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe21[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe21[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe21[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe21[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe21[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe21[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe21[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),	
	.dout_w_b1_30(dout_w_b1_pe21[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe21[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe21[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe21[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe21[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe21[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe21[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe21[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe21[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe21[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[9]),
	.dout_psum0_00(psum0_pe21[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe21[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe21[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe21[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe21[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe21[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe21[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe21[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe21[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe21[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe21[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe21[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe21[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe21[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe21[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe21[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe21[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe21[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe21[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe21[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe21[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe21[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe21[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe21[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe21[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[9]),
	.dout_psum1_00(psum1_pe21[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe21[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe21[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe21[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe21[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe21[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe21[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe21[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe21[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe21[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe21[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe21[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe21[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe21[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe21[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe21[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe21[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe21[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe21[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe21[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe21[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe21[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe21[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe21[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe21[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_norm#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_22(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe21),
	.din_fm_00(dout_fm_pe21[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe21[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe21[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe21[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe21[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe21[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe21[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe21[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe21[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe21[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe21[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe21[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe21[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe21[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(dout_fm_pe21[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(dout_fm_pe21[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe21[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_fm_32(dout_fm_pe21[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe21[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe21[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe21[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe21[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe21[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe21[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe21[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe12),
	.din_w_b0_00(dout_w_b0_pe12[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe12[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe12[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe12[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe12[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe12[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe12[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe12[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe12[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe12[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe12[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe12[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe12[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe12[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe12[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe12[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe12[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe12[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe12[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe12[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe12[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe12[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe12[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe12[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe12[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe12),
	.din_w_b1_00(dout_w_b1_pe12[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe12[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe12[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe12[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe12[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe12[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe12[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe12[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe12[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe12[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe12[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe12[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe12[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe12[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe12[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe12[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe12[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe12[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe12[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe12[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe12[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe12[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe12[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe12[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe12[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe22),
	.dout_fm_00(dout_fm_pe22[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe22[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe22[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe22[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe22[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe22[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe22[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe22[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe22[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe22[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe22[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe22[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe22[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe22[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe22[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe22[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe22[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe22[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe22[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe22[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe22[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe22[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe22[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe22[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe22[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe22),
	.dout_w_b0_00(dout_w_b0_pe22[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe22[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe22[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe22[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b0_04(dout_w_b0_pe22[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe22[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe22[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe22[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe22[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe22[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe22[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe22[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe22[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe22[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe22[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe22[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe22[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe22[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe22[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe22[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe22[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe22[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe22[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe22[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),	
	.dout_w_b0_44(dout_w_b0_pe22[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk	
	.en_out_w_b1(en_out_w_b1_pe22),
	.dout_w_b1_00(dout_w_b1_pe22[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe22[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe22[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe22[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b1_04(dout_w_b1_pe22[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe22[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe22[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe22[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe22[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe22[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe22[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe22[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe22[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe22[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe22[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),	
	.dout_w_b1_30(dout_w_b1_pe22[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe22[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe22[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe22[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe22[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe22[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe22[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe22[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe22[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe22[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[10]),
	.dout_psum0_00(psum0_pe22[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe22[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe22[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe22[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe22[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe22[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe22[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe22[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe22[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe22[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe22[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe22[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe22[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe22[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe22[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe22[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe22[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe22[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe22[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe22[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe22[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe22[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe22[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe22[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe22[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[10]),
	.dout_psum1_00(psum1_pe22[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe22[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe22[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe22[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe22[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe22[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe22[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe22[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe22[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe22[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe22[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe22[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe22[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe22[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe22[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe22[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe22[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe22[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe22[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe22[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe22[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe22[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe22[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe22[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe22[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_right#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_23(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe22),
	.din_fm_00(dout_fm_pe22[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe22[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe22[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe22[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe22[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe22[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe22[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe22[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe22[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe22[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe22[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe22[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe22[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe22[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(dout_fm_pe22[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(dout_fm_pe22[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe22[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_fm_32(dout_fm_pe22[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe22[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe22[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe22[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe22[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe22[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe22[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe22[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe13),
	.din_w_b0_00(dout_w_b0_pe13[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe13[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe13[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe13[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe13[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe13[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe13[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe13[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe13[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe13[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe13[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe13[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe13[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe13[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe13[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe13[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe13[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe13[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe13[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe13[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe13[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe13[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe13[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe13[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe13[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe13),
	.din_w_b1_00(dout_w_b1_pe13[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe13[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe13[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe13[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe13[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe13[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe13[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe13[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe13[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe13[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe13[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe13[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe13[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe13[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe13[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe13[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe13[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe13[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe13[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe13[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe13[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe13[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe13[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe13[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe13[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0 delay 1 clk
	.en_out_w_b0(en_out_w_b0_pe23),
	.dout_w_b0_00(dout_w_b0_pe23[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b0_01(dout_w_b0_pe23[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b0_02(dout_w_b0_pe23[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b0_03(dout_w_b0_pe23[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b0_04(dout_w_b0_pe23[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b0_10(dout_w_b0_pe23[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b0_11(dout_w_b0_pe23[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b0_12(dout_w_b0_pe23[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b0_13(dout_w_b0_pe23[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b0_14(dout_w_b0_pe23[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b0_20(dout_w_b0_pe23[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b0_21(dout_w_b0_pe23[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b0_22(dout_w_b0_pe23[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b0_23(dout_w_b0_pe23[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b0_24(dout_w_b0_pe23[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_w_b0_30(dout_w_b0_pe23[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b0_31(dout_w_b0_pe23[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b0_32(dout_w_b0_pe23[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b0_33(dout_w_b0_pe23[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b0_34(dout_w_b0_pe23[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b0_40(dout_w_b0_pe23[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b0_41(dout_w_b0_pe23[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b0_42(dout_w_b0_pe23[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b0_43(dout_w_b0_pe23[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),	
	.dout_w_b0_44(dout_w_b0_pe23[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1 delay 1 clk	
	.en_out_w_b1(en_out_w_b1_pe23),
	.dout_w_b1_00(dout_w_b1_pe23[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_w_b1_01(dout_w_b1_pe23[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_w_b1_02(dout_w_b1_pe23[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_w_b1_03(dout_w_b1_pe23[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),	
	.dout_w_b1_04(dout_w_b1_pe23[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_w_b1_10(dout_w_b1_pe23[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_w_b1_11(dout_w_b1_pe23[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_w_b1_12(dout_w_b1_pe23[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_w_b1_13(dout_w_b1_pe23[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_w_b1_14(dout_w_b1_pe23[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_w_b1_20(dout_w_b1_pe23[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_w_b1_21(dout_w_b1_pe23[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_w_b1_22(dout_w_b1_pe23[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_w_b1_23(dout_w_b1_pe23[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_w_b1_24(dout_w_b1_pe23[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),	
	.dout_w_b1_30(dout_w_b1_pe23[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_w_b1_31(dout_w_b1_pe23[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_w_b1_32(dout_w_b1_pe23[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_w_b1_33(dout_w_b1_pe23[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_w_b1_34(dout_w_b1_pe23[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_w_b1_40(dout_w_b1_pe23[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_w_b1_41(dout_w_b1_pe23[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_w_b1_42(dout_w_b1_pe23[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_w_b1_43(dout_w_b1_pe23[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_w_b1_44(dout_w_b1_pe23[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[11]),
	.dout_psum0_00(psum0_pe23[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe23[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe23[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe23[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe23[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe23[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe23[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe23[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe23[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe23[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe23[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe23[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe23[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe23[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe23[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe23[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe23[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe23[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe23[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe23[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe23[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe23[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe23[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe23[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe23[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[11]),
	.dout_psum1_00(psum1_pe23[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe23[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe23[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe23[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe23[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe23[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe23[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe23[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe23[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe23[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe23[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe23[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe23[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe23[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe23[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe23[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe23[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe23[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe23[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe23[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe23[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe23[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe23[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe23[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe23[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);


pe_bottom#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_30(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_fm[3]),
	.din_fm_00(din_fm_c3[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(din_fm_c3[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(din_fm_c3[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(din_fm_c3[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(din_fm_c3[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(din_fm_c3[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(din_fm_c3[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(din_fm_c3[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(din_fm_c3[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(din_fm_c3[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(din_fm_c3[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(din_fm_c3[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(din_fm_c3[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(din_fm_c3[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(din_fm_c3[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(din_fm_c3[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(din_fm_c3[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_fm_32(din_fm_c3[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(din_fm_c3[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(din_fm_c3[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(din_fm_c3[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(din_fm_c3[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(din_fm_c3[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(din_fm_c3[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(din_fm_c3[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe20),
	.din_w_b0_00(dout_w_b0_pe20[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe20[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe20[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe20[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe20[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe20[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe20[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe20[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe20[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe20[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe20[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe20[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe20[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe20[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe20[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe20[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe20[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe20[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe20[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe20[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe20[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe20[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe20[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe20[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe20[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe20), // ok
	.din_w_b1_00(dout_w_b1_pe20[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe20[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe20[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe20[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe20[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe20[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe20[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe20[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe20[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe20[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe20[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe20[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe20[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe20[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe20[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe20[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe20[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe20[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe20[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe20[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe20[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe20[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe20[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe20[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe20[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe30),
	.dout_fm_00(dout_fm_pe30[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe30[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe30[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe30[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe30[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe30[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe30[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe30[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe30[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe30[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe30[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe30[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe30[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe30[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe30[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe30[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe30[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe30[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe30[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe30[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe30[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe30[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe30[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe30[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe30[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[12]),
	.dout_psum0_00(psum0_pe30[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe30[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe30[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe30[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe30[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe30[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe30[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe30[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe30[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe30[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe30[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe30[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe30[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe30[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe30[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe30[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe30[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe30[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe30[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe30[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe30[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe30[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe30[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe30[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe30[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[12]),
	.dout_psum1_00(psum1_pe30[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe30[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe30[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe30[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe30[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe30[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe30[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe30[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe30[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe30[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe30[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe30[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe30[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe30[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe30[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe30[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe30[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe30[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe30[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe30[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe30[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe30[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe30[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe30[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe30[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_bottom#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_31(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe30),
	.din_fm_00(dout_fm_pe30[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe30[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe30[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe30[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe30[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe30[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe30[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe30[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe30[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe30[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe30[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe30[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe30[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe30[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(dout_fm_pe30[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(dout_fm_pe30[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe30[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_fm_32(dout_fm_pe30[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe30[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe30[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe30[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe30[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe30[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe30[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe30[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe21),
	.din_w_b0_00(dout_w_b0_pe21[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe21[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe21[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe21[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe21[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe21[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe21[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe21[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe21[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe21[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe21[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe21[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe21[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe21[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe21[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe21[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe21[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe21[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe21[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe21[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe21[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe21[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe21[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe21[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe21[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe21),
	.din_w_b1_00(dout_w_b1_pe21[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe21[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe21[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe21[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe21[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe21[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe21[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe21[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe21[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe21[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe21[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe21[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe21[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe21[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe21[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe21[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe21[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe21[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe21[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe21[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe21[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe21[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe21[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe21[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe21[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe31),
	.dout_fm_00(dout_fm_pe31[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe31[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe31[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe31[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe31[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe31[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe31[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe31[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe31[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe31[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe31[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe31[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe31[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe31[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe31[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe31[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe31[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe31[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe31[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe31[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe31[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe31[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe31[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe31[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe31[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[13]),
	.dout_psum0_00(psum0_pe31[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe31[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe31[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe31[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe31[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe31[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe31[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe31[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe31[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe31[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe31[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe31[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe31[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe31[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe31[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe31[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe31[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe31[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe31[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe31[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe31[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe31[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe31[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe31[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe31[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[13]),
	.dout_psum1_00(psum1_pe31[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe31[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe31[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe31[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe31[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe31[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe31[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe31[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe31[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe31[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe31[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe31[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe31[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe31[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe31[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe31[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe31[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe31[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe31[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe31[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe31[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe31[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe31[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe31[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe31[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_bottom#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_32(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe31),
	.din_fm_00(dout_fm_pe31[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe31[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe31[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe31[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe31[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe31[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe31[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe31[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe31[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe31[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe31[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe31[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe31[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe31[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(dout_fm_pe31[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(dout_fm_pe31[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe31[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_fm_32(dout_fm_pe31[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe31[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe31[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe31[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe31[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe31[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe31[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe31[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe22),
	.din_w_b0_00(dout_w_b0_pe22[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe22[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe22[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe22[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe22[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe22[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe22[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe22[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe22[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe22[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe22[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe22[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe22[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe22[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe22[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe22[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe22[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe22[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe22[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe22[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe22[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe22[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe22[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe22[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe22[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe22),
	.din_w_b1_00(dout_w_b1_pe22[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe22[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe22[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe22[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe22[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe22[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe22[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe22[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe22[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe22[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe22[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe22[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe22[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe22[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe22[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe22[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe22[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe22[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe22[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe22[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe22[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe22[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe22[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe22[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe22[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input feature map delay 1 clk
	.en_out_fm(en_out_fm_pe32),
	.dout_fm_00(dout_fm_pe32[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.dout_fm_01(dout_fm_pe32[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.dout_fm_02(dout_fm_pe32[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.dout_fm_03(dout_fm_pe32[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.dout_fm_04(dout_fm_pe32[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.dout_fm_10(dout_fm_pe32[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.dout_fm_11(dout_fm_pe32[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.dout_fm_12(dout_fm_pe32[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.dout_fm_13(dout_fm_pe32[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.dout_fm_14(dout_fm_pe32[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.dout_fm_20(dout_fm_pe32[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.dout_fm_21(dout_fm_pe32[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.dout_fm_22(dout_fm_pe32[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.dout_fm_23(dout_fm_pe32[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.dout_fm_24(dout_fm_pe32[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.dout_fm_30(dout_fm_pe32[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.dout_fm_31(dout_fm_pe32[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.dout_fm_32(dout_fm_pe32[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.dout_fm_33(dout_fm_pe32[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.dout_fm_34(dout_fm_pe32[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.dout_fm_40(dout_fm_pe32[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.dout_fm_41(dout_fm_pe32[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.dout_fm_42(dout_fm_pe32[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.dout_fm_43(dout_fm_pe32[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.dout_fm_44(dout_fm_pe32[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[14]),
	.dout_psum0_00(psum0_pe32[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe32[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe32[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe32[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe32[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe32[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe32[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe32[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe32[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe32[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe32[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe32[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe32[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe32[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe32[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe32[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe32[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe32[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe32[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe32[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe32[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe32[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe32[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe32[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe32[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[14]),
	.dout_psum1_00(psum1_pe32[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe32[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe32[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe32[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe32[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe32[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe32[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe32[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe32[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe32[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe32[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe32[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe32[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe32[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe32[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe32[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe32[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe32[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe32[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe32[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe32[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe32[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe32[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe32[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe32[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

pe_lrcorner#(
	.DATA_WIDTH_I(DATA_WIDTH_I),
	.DATA_WIDTH_O(DATA_WIDTH_O)
) pe_33(
	.clk(clk),
	.rst(rst_d1),
	// input feature map
	.en_fm(en_out_fm_pe32),
	.din_fm_00(dout_fm_pe32[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_fm_01(dout_fm_pe32[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_fm_02(dout_fm_pe32[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_fm_03(dout_fm_pe32[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_fm_04(dout_fm_pe32[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_fm_10(dout_fm_pe32[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_fm_11(dout_fm_pe32[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_fm_12(dout_fm_pe32[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_fm_13(dout_fm_pe32[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_fm_14(dout_fm_pe32[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_fm_20(dout_fm_pe32[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_fm_21(dout_fm_pe32[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_fm_22(dout_fm_pe32[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_fm_23(dout_fm_pe32[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_fm_24(dout_fm_pe32[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_fm_30(dout_fm_pe32[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_fm_31(dout_fm_pe32[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_fm_32(dout_fm_pe32[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_fm_33(dout_fm_pe32[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_fm_34(dout_fm_pe32[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_fm_40(dout_fm_pe32[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_fm_41(dout_fm_pe32[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_fm_42(dout_fm_pe32[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_fm_43(dout_fm_pe32[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_fm_44(dout_fm_pe32[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 0
	.en_w_b0(en_out_w_b0_pe23),
	.din_w_b0_00(dout_w_b0_pe23[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b0_01(dout_w_b0_pe23[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b0_02(dout_w_b0_pe23[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b0_03(dout_w_b0_pe23[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b0_04(dout_w_b0_pe23[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b0_10(dout_w_b0_pe23[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b0_11(dout_w_b0_pe23[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b0_12(dout_w_b0_pe23[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b0_13(dout_w_b0_pe23[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b0_14(dout_w_b0_pe23[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b0_20(dout_w_b0_pe23[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b0_21(dout_w_b0_pe23[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b0_22(dout_w_b0_pe23[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b0_23(dout_w_b0_pe23[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b0_24(dout_w_b0_pe23[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b0_30(dout_w_b0_pe23[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b0_31(dout_w_b0_pe23[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),	
	.din_w_b0_32(dout_w_b0_pe23[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b0_33(dout_w_b0_pe23[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b0_34(dout_w_b0_pe23[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b0_40(dout_w_b0_pe23[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b0_41(dout_w_b0_pe23[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b0_42(dout_w_b0_pe23[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b0_43(dout_w_b0_pe23[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b0_44(dout_w_b0_pe23[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// input weight batch 1
	.en_w_b1(en_out_w_b1_pe23),
	.din_w_b1_00(dout_w_b1_pe23[DATA_WIDTH_I*1-1 :DATA_WIDTH_I*0 ]),.din_w_b1_01(dout_w_b1_pe23[DATA_WIDTH_I*2-1 :DATA_WIDTH_I*1 ]),
	.din_w_b1_02(dout_w_b1_pe23[DATA_WIDTH_I*3-1 :DATA_WIDTH_I*2 ]),.din_w_b1_03(dout_w_b1_pe23[DATA_WIDTH_I*4-1 :DATA_WIDTH_I*3 ]),
	.din_w_b1_04(dout_w_b1_pe23[DATA_WIDTH_I*5-1 :DATA_WIDTH_I*4 ]),
	.din_w_b1_10(dout_w_b1_pe23[DATA_WIDTH_I*6-1 :DATA_WIDTH_I*5 ]),.din_w_b1_11(dout_w_b1_pe23[DATA_WIDTH_I*7-1 :DATA_WIDTH_I*6 ]),
	.din_w_b1_12(dout_w_b1_pe23[DATA_WIDTH_I*8-1 :DATA_WIDTH_I*7 ]),.din_w_b1_13(dout_w_b1_pe23[DATA_WIDTH_I*9-1 :DATA_WIDTH_I*8 ]),
	.din_w_b1_14(dout_w_b1_pe23[DATA_WIDTH_I*10-1:DATA_WIDTH_I*9 ]),
	.din_w_b1_20(dout_w_b1_pe23[DATA_WIDTH_I*11-1:DATA_WIDTH_I*10]),.din_w_b1_21(dout_w_b1_pe23[DATA_WIDTH_I*12-1:DATA_WIDTH_I*11]),
	.din_w_b1_22(dout_w_b1_pe23[DATA_WIDTH_I*13-1:DATA_WIDTH_I*12]),.din_w_b1_23(dout_w_b1_pe23[DATA_WIDTH_I*14-1:DATA_WIDTH_I*13]),
	.din_w_b1_24(dout_w_b1_pe23[DATA_WIDTH_I*15-1:DATA_WIDTH_I*14]),
	.din_w_b1_30(dout_w_b1_pe23[DATA_WIDTH_I*16-1:DATA_WIDTH_I*15]),.din_w_b1_31(dout_w_b1_pe23[DATA_WIDTH_I*17-1:DATA_WIDTH_I*16]),
	.din_w_b1_32(dout_w_b1_pe23[DATA_WIDTH_I*18-1:DATA_WIDTH_I*17]),.din_w_b1_33(dout_w_b1_pe23[DATA_WIDTH_I*19-1:DATA_WIDTH_I*18]),
	.din_w_b1_34(dout_w_b1_pe23[DATA_WIDTH_I*20-1:DATA_WIDTH_I*19]),
	.din_w_b1_40(dout_w_b1_pe23[DATA_WIDTH_I*21-1:DATA_WIDTH_I*20]),.din_w_b1_41(dout_w_b1_pe23[DATA_WIDTH_I*22-1:DATA_WIDTH_I*21]),
	.din_w_b1_42(dout_w_b1_pe23[DATA_WIDTH_I*23-1:DATA_WIDTH_I*22]),.din_w_b1_43(dout_w_b1_pe23[DATA_WIDTH_I*24-1:DATA_WIDTH_I*23]),
	.din_w_b1_44(dout_w_b1_pe23[DATA_WIDTH_I*25-1:DATA_WIDTH_I*24]),
	// output partial sum 0	
	.en_psum0(en_psum0[15]),
	.dout_psum0_00(psum0_pe33[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum0_01(psum0_pe33[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum0_02(psum0_pe33[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum0_03(psum0_pe33[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum0_04(psum0_pe33[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum0_10(psum0_pe33[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum0_11(psum0_pe33[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum0_12(psum0_pe33[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum0_13(psum0_pe33[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum0_14(psum0_pe33[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),	
	.dout_psum0_20(psum0_pe33[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum0_21(psum0_pe33[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),	
	.dout_psum0_22(psum0_pe33[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum0_23(psum0_pe33[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum0_24(psum0_pe33[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum0_30(psum0_pe33[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum0_31(psum0_pe33[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum0_32(psum0_pe33[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum0_33(psum0_pe33[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum0_34(psum0_pe33[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum0_40(psum0_pe33[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum0_41(psum0_pe33[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum0_42(psum0_pe33[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum0_43(psum0_pe33[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum0_44(psum0_pe33[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24]),
	// output partial sum 1	
	.en_psum1(en_psum1[15]),
	.dout_psum1_00(psum1_pe33[DATA_WIDTH_O*1-1 :DATA_WIDTH_O*0 ]),.dout_psum1_01(psum1_pe33[DATA_WIDTH_O*2-1 :DATA_WIDTH_O*1 ]),
	.dout_psum1_02(psum1_pe33[DATA_WIDTH_O*3-1 :DATA_WIDTH_O*2 ]),.dout_psum1_03(psum1_pe33[DATA_WIDTH_O*4-1 :DATA_WIDTH_O*3 ]),
	.dout_psum1_04(psum1_pe33[DATA_WIDTH_O*5-1 :DATA_WIDTH_O*4 ]),
	.dout_psum1_10(psum1_pe33[DATA_WIDTH_O*6-1 :DATA_WIDTH_O*5 ]),.dout_psum1_11(psum1_pe33[DATA_WIDTH_O*7-1 :DATA_WIDTH_O*6 ]),
	.dout_psum1_12(psum1_pe33[DATA_WIDTH_O*8-1 :DATA_WIDTH_O*7 ]),.dout_psum1_13(psum1_pe33[DATA_WIDTH_O*9-1 :DATA_WIDTH_O*8 ]),
	.dout_psum1_14(psum1_pe33[DATA_WIDTH_O*10-1:DATA_WIDTH_O*9 ]),
	.dout_psum1_20(psum1_pe33[DATA_WIDTH_O*11-1:DATA_WIDTH_O*10]),.dout_psum1_21(psum1_pe33[DATA_WIDTH_O*12-1:DATA_WIDTH_O*11]),
	.dout_psum1_22(psum1_pe33[DATA_WIDTH_O*13-1:DATA_WIDTH_O*12]),.dout_psum1_23(psum1_pe33[DATA_WIDTH_O*14-1:DATA_WIDTH_O*13]),
	.dout_psum1_24(psum1_pe33[DATA_WIDTH_O*15-1:DATA_WIDTH_O*14]),	
	.dout_psum1_30(psum1_pe33[DATA_WIDTH_O*16-1:DATA_WIDTH_O*15]),.dout_psum1_31(psum1_pe33[DATA_WIDTH_O*17-1:DATA_WIDTH_O*16]),
	.dout_psum1_32(psum1_pe33[DATA_WIDTH_O*18-1:DATA_WIDTH_O*17]),.dout_psum1_33(psum1_pe33[DATA_WIDTH_O*19-1:DATA_WIDTH_O*18]),
	.dout_psum1_34(psum1_pe33[DATA_WIDTH_O*20-1:DATA_WIDTH_O*19]),	
	.dout_psum1_40(psum1_pe33[DATA_WIDTH_O*21-1:DATA_WIDTH_O*20]),.dout_psum1_41(psum1_pe33[DATA_WIDTH_O*22-1:DATA_WIDTH_O*21]),
	.dout_psum1_42(psum1_pe33[DATA_WIDTH_O*23-1:DATA_WIDTH_O*22]),.dout_psum1_43(psum1_pe33[DATA_WIDTH_O*24-1:DATA_WIDTH_O*23]),
	.dout_psum1_44(psum1_pe33[DATA_WIDTH_O*25-1:DATA_WIDTH_O*24])
);

endmodule

